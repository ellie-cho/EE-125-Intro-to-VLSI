library ieee;
use ieee.std_logic_1164.all;

entity vga is
	 generic (
	 H_LOW: natural := 96;
	 HBP: natural := 48;
	 H_HIGH: natural := 640;
	 HFP: natural := 16;
	 V_LOW: natural := 2;
	 VBP: natural := 33;
	 V_HIGH: natural := 480;
	 VFP: natural := 10);
	 port (
	 clk: in std_logic; --50MHz system clock
	 R_switch, G_switch, B_switch: in std_logic;
	 Hsync, Vsync: out std_logic;
	 R, G, B: out std_logic_vector(3 downto 0);
	 BLANKn, SYNCn : out std_logic);
	 
end entity;

architecture rtl of vga is
	 signal Hactive, Vactive, dena: std_logic;
	 signal clk_vga, Hsyn, Vsyn: std_logic;
	 type rgb_array is array (1 to 48) of std_logic_vector(3 downto 0);
	 type img_array is array (1 to 48) of rgb_array;
    constant r_image_data : img_array := 
	 (("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0110", "1000", "0100", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0010", "0101", "0111", "1001", "1010", "1010", "0101", "0000", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0010", "0101", "1000", "1001", "1010", "1010", "1010", "1010", "1010", "1000", "0010", "0100", "0100", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0010", "0110", "1000", "1010", "1010", "1010", "1010", "1010", "1001", "1010", "1000", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "0110", "0100", "0100", "0010", "0010", "0010", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0100", "0111", "1000", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1000", "1010", "0011", "0100", "0011", "0011", "0011", "0100", "0100", "0101", "0101", "0110", "0111", "0111", "1000", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "0101", "0010", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0010", "0100", "0111", "1000", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1000", "1001", "0011", "0100", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0100", "0100", "0100", "0100", "0111", "1001", "0111", "0100", "0101", "0110", "1010", "0010", "0010", "0011", "0011"), ("0011", "0011", "0011", "0010", "0110", "0111", "1000", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1000", "1000", "0011", "0100", "0011", "0010", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0100", "0100", "0111", "1010", "1001", "0100", "0101", "0101", "1010", "0001", "0010", "0011", "0011"), ("0011", "0011", "0011", "0100", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "0111", "0111", "0011", "0011", "0011", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0011", "0100", "0101", "1010", "1010", "0011", "0100", "0100", "1010", "0000", "0010", "0011", "0011"), ("0011", "0011", "1001", "0101", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "0111", "0111", "0010", "0011", "0011", "0001", "0001", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0100", "1010", "1010", "0011", "0100", "0100", "1010", "0100", "1001", "0011", "0011"), ("0011", "1001", "1000", "0111", "1000", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1000", "1000", "0111", "0110", "0010", "0010", "0010", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0010", "0011", "0100", "1010", "1010", "0010", "0100", "0011", "1001", "0111", "1001", "1001", "0011"), ("1001", "1000", "0010", "0001", "0010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1010", "1000", "1000", "1000", "1000", "0111", "0101", "0101", "0111", "0101", "0010", "0010", "0010", "0001", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0011", "1001", "1010", "0010", "0011", "0100", "1000", "0001", "0011", "1000", "1001"), ("1001", "1000", "0001", "0000", "0000", "0111", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "0111", "0110", "0110", "0101", "0101", "0101", "0011", "0010", "0110", "0100", "0010", "0010", "0010", "0001", "0000", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0001", "0010", "0111", "1001", "0001", "0010", "0011", "0110", "0000", "0001", "1000", "1001"), ("1001", "1000", "0001", "0000", "0000", "0100", "0111", "0110", "0111", "0110", "0101", "0101", "0100", "0100", "0011", "0100", "0001", "0001", "0011", "0001", "0000", "0101", "0011", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0101", "0111", "0001", "0010", "0011", "0101", "0000", "0010", "1000", "1001"), ("1001", "1000", "0110", "0110", "0110", "0111", "1000", "0111", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0111", "0111", "0110", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0111", "0110", "0110", "0110", "0111", "1000", "1000", "0110", "0111", "0111", "0111", "0110", "0111", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1000", "1000", "1000", "1000", "1001", "1001", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1001", "1000", "0111", "0101", "0100", "0011", "0011", "0100", "0101", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1001", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1000", "0111", "0100", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0010", "0100", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1001", "0111", "1000", "1001"), ("1001", "1000", "0111", "0111", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1000", "0101", "0010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0110", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "0110", "1000", "1001"), ("1001", "1000", "0111", "0110", "0111", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0110", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "1000", "1001"), ("1001", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "0111", "0110", "0010", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0100", "0100", "0011", "0001", "0000", "0000", "0001", "0011", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "1001"), ("1001", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1000", "0011", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0010", "0011", "0100", "0100", "0100", "0001", "0000", "0000", "0010", "0100", "1000", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "1001"), ("1001", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "0110", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0011", "0011", "0001", "0001", "0000", "0000", "0010", "0111", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1000", "0100", "0001", "0000", "0000", "0010", "0001", "0001", "0001", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "0101", "1000", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0011", "0001", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0011", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0000", "0000", "0001", "0001", "0010", "0001", "0000", "0000", "0001", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "1001"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0000", "0000", "0001", "0001", "0010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0001", "0001", "0000", "0000", "0010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "1001"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0001", "0000", "0001", "0001", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0001", "0001", "0000", "0000", "0011", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1001", "0100", "0001", "0000", "0001", "0001", "0010", "0011", "0001", "0000", "0000", "0000", "0000", "0001", "0011", "0001", "0001", "0000", "0000", "0000", "0101", "1001", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1001", "0111", "0001", "0000", "0000", "0001", "0001", "0010", "0011", "0010", "0001", "0001", "0010", "0011", "0010", "0001", "0001", "0000", "0000", "0000", "1000", "1001", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1010", "0011", "0000", "0000", "0001", "0001", "0001", "0010", "0010", "0011", "0011", "0010", "0010", "0001", "0001", "0000", "0000", "0000", "0011", "1010", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1001", "0111", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "1000", "1001", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "1001", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1010", "0101", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0001", "0110", "1010", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1001", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1010", "0101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0101", "1010", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0111", "1000"), ("1000", "0111", "0111", "0110", "0110", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1010", "0111", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0111", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0110", "0111", "1000", "1000"), ("1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1010", "1010", "0111", "0100", "0010", "0001", "0001", "0010", "0100", "0111", "1010", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1001", "1001", "1001", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001"), ("0011", "0011", "0011", "0011", "0010", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0110", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0110", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0010", "0010", "0011", "0011", "0011"), ("0011", "0011", "0011", "0000", "0001", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0101", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0001", "0000", "0011", "0011", "0011"), ("0011", "0011", "0010", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0000", "0000", "0010", "0011", "0011", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0011", "0011", "0010", "0000", "0000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0010", "0011", "0011"), ("0011", "0011", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0011", "0011"), ("0011", "0011", "0011", "0010", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0000", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0010", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"));	 
	 constant g_image_data: img_array := 
	(("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "0110", "1000", "0100", "0010", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "0010", "0101", "0111", "1001", "1010", "1010", "0101", "0000", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "0010", "0101", "1000", "1001", "1010", "1010", "1010", "1001", "1001", "1000", "0010", "0100", "0100", "0010", "0010", "0010", "0010", "0010", "0010", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "0010", "0110", "1000", "1010", "1010", "1010", "1001", "1001", "1000", "1010", "1000", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "0110", "0100", "0100", "0010", "0010", "0010", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "0100", "0111", "1000", "1010", "1010", "1010", "1001", "1001", "1001", "1010", "1001", "1000", "1010", "0011", "0100", "0011", "0010", "0011", "0100", "0100", "0101", "0101", "0110", "0111", "0111", "1000", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "0101", "0010", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0010", "0100", "0111", "1000", "1010", "1010", "1010", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1001", "0111", "1001", "0011", "0100", "0011", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0100", "0100", "0111", "1001", "0111", "0100", "0101", "0110", "1010", "0010", "0010", "0100", "0100"), ("0100", "0100", "0100", "0010", "0110", "0111", "1000", "1010", "1010", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "0111", "1000", "0010", "0011", "0011", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0011", "0011", "0100", "0110", "1010", "1001", "0100", "0101", "0101", "1010", "0001", "0010", "0100", "0100"), ("0100", "0100", "0100", "0100", "1010", "1010", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "0111", "0111", "0010", "0011", "0010", "0001", "0001", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0101", "1010", "1001", "0011", "0100", "0011", "1010", "0000", "0010", "0100", "0100"), ("0100", "0100", "1001", "0101", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0111", "0111", "0010", "0010", "0010", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0010", "0011", "0100", "1010", "1010", "0010", "0100", "0011", "1001", "0100", "1001", "0100", "0100"), ("0100", "1001", "1000", "0111", "1000", "1010", "1010", "1010", "1010", "1001", "1010", "1001", "1001", "1001", "1000", "1001", "1000", "1000", "1000", "0111", "0110", "0110", "0110", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0100", "1010", "1010", "0010", "0011", "0011", "1001", "0111", "1000", "1001", "0100"), ("1001", "1000", "0010", "0001", "0010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0111", "0111", "0110", "0111", "0101", "0100", "0011", "0110", "0101", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "1001", "1010", "0001", "0011", "0011", "1000", "0001", "0011", "1000", "1001"), ("1001", "1000", "0001", "0000", "0000", "0111", "1000", "1000", "1000", "1000", "1000", "0110", "0110", "0101", "0101", "0101", "0011", "0100", "0100", "0010", "0001", "0110", "0100", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0111", "1001", "0000", "0010", "0011", "0110", "0000", "0001", "1000", "1001"), ("1001", "1000", "0001", "0000", "0000", "0100", "0111", "0101", "0110", "0101", "0100", "0011", "0010", "0011", "0010", "0011", "0001", "0001", "0010", "0000", "0000", "0101", "0010", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0101", "0111", "0000", "0010", "0011", "0101", "0000", "0010", "1000", "1001"), ("1001", "1000", "0110", "0110", "0110", "0111", "1000", "0111", "0111", "0111", "0111", "0111", "0110", "0111", "0110", "0110", "0110", "0110", "0111", "0110", "0110", "1000", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "1000", "0110", "0111", "0111", "0111", "0110", "0111", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1001", "1000", "0111", "0101", "0100", "0011", "0011", "0100", "0101", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1001", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1000", "0111", "0011", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0010", "0100", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1001", "0111", "1000", "1001"), ("1001", "1000", "0111", "0111", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0101", "0010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0110", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "0110", "1000", "1001"), ("1001", "1000", "0111", "0110", "0111", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0110", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "1000", "1001"), ("1001", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "0111", "0110", "0010", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0100", "0100", "0011", "0001", "0000", "0000", "0001", "0011", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "1001"), ("1001", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1000", "0011", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0010", "0011", "0100", "0100", "0100", "0001", "0000", "0000", "0010", "0100", "1000", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "1001"), ("1001", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "0110", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0011", "0011", "0001", "0001", "0000", "0000", "0010", "0111", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1000", "0100", "0001", "0000", "0000", "0010", "0001", "0001", "0001", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "0101", "1000", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0011", "0001", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0011", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0000", "0000", "0001", "0001", "0010", "0001", "0000", "0000", "0001", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "1001"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0000", "0000", "0001", "0001", "0010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0001", "0001", "0000", "0000", "0010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "1001"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0001", "0000", "0001", "0001", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0001", "0001", "0000", "0000", "0011", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1001", "0100", "0001", "0000", "0001", "0001", "0010", "0011", "0001", "0000", "0000", "0000", "0000", "0001", "0011", "0001", "0001", "0000", "0000", "0000", "0101", "1001", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1001", "0111", "0001", "0000", "0000", "0001", "0001", "0010", "0011", "0010", "0001", "0001", "0010", "0011", "0010", "0001", "0001", "0000", "0000", "0000", "1000", "1001", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1010", "0011", "0000", "0000", "0001", "0001", "0001", "0010", "0010", "0011", "0011", "0010", "0010", "0001", "0001", "0000", "0000", "0000", "0011", "1010", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1001", "0111", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "1000", "1001", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "1001", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1010", "0101", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0001", "0110", "1010", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1001", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1010", "0101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0101", "1010", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0111", "1000"), ("1000", "0111", "0111", "0110", "0110", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1010", "0111", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0111", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0110", "0111", "1000", "1000"), ("1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1010", "1010", "0111", "0100", "0010", "0001", "0001", "0010", "0100", "0111", "1010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1001", "1001", "1001", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001"), ("0100", "0100", "0100", "0011", "0010", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0110", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0110", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0010", "0010", "0100", "0100", "0100"), ("0100", "0100", "0100", "0000", "0001", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0101", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0001", "0000", "0100", "0100", "0100"), ("0100", "0100", "0010", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0000", "0000", "0010", "0011", "0011", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0011", "0011", "0010", "0000", "0000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0010", "0100", "0100"), ("0100", "0100", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0100", "0100"), ("0100", "0100", "0100", "0010", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0000", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0010", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"), ("0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100"));	 
	 constant b_image_data: img_array := 
	 (("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0110", "1000", "0100", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0010", "0101", "0111", "1001", "1010", "1010", "0101", "0000", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0010", "0101", "1000", "1001", "1010", "1001", "1010", "1001", "1000", "1000", "0010", "0100", "0100", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0010", "0110", "1000", "1010", "1010", "1001", "1001", "1000", "0111", "1010", "1000", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "0110", "0100", "0100", "0010", "0010", "0010", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0100", "0111", "1000", "1010", "1010", "1001", "1001", "1000", "1001", "1001", "1001", "0111", "1010", "0011", "0100", "0011", "0010", "0011", "0100", "0100", "0101", "0101", "0110", "0111", "0111", "1000", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "0101", "0010", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0010", "0100", "0111", "1000", "1010", "1010", "1001", "1001", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "0111", "1001", "0011", "0100", "0011", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0100", "0100", "0110", "1001", "0111", "0100", "0101", "0110", "1010", "0010", "0010", "0011", "0011"), ("0011", "0011", "0011", "0010", "0110", "0111", "1000", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0111", "1000", "0010", "0011", "0011", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0011", "0011", "0100", "0110", "1010", "1001", "0100", "0101", "0101", "1010", "0001", "0010", "0011", "0011"), ("0011", "0011", "0011", "0100", "1010", "1010", "1001", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "0111", "0111", "0010", "0011", "0010", "0001", "0001", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0011", "0011", "0101", "1010", "1001", "0011", "0100", "0011", "1010", "0000", "0010", "0011", "0011"), ("0011", "0011", "1001", "0101", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0110", "0111", "0010", "0010", "0010", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0010", "0011", "0100", "1010", "1010", "0010", "0100", "0011", "1001", "0100", "1001", "0011", "0011"), ("0011", "1001", "1000", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "0111", "1000", "0111", "0111", "0111", "0101", "0101", "0110", "0110", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0100", "1010", "1010", "0010", "0011", "0011", "1001", "0111", "1001", "1001", "0011"), ("1001", "1000", "0010", "0001", "0010", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0101", "0101", "0101", "0101", "0100", "0010", "0010", "0110", "0101", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "1001", "1001", "0001", "0011", "0011", "1000", "0001", "0011", "1000", "1001"), ("1001", "1000", "0001", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0101", "0101", "0100", "0100", "0100", "0010", "0010", "0010", "0001", "0000", "0110", "0100", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0111", "1001", "0000", "0010", "0011", "0110", "0000", "0001", "1000", "1001"), ("1001", "1000", "0001", "0000", "0000", "0100", "0110", "0011", "0101", "0100", "0010", "0010", "0001", "0010", "0001", "0010", "0000", "0000", "0001", "0000", "0000", "0101", "0010", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0101", "0111", "0000", "0010", "0011", "0101", "0000", "0010", "1000", "1001"), ("1001", "1000", "0110", "0110", "0110", "0111", "1000", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "1000", "0110", "0111", "0111", "1000", "0110", "0111", "1000", "1001"), ("1001", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1001", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1001", "1000", "0111", "0101", "0100", "0011", "0011", "0100", "0101", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1001", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1000", "0111", "0011", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0010", "0100", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1001", "0111", "1000", "1001"), ("1001", "1000", "0111", "0111", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0101", "0010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0110", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "0110", "1000", "1001"), ("1001", "1000", "0111", "0110", "0111", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "0101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0110", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "1000", "1000", "1001"), ("1001", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "0111", "0110", "0010", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0100", "0100", "0011", "0001", "0000", "0000", "0001", "0011", "0110", "0111", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "1001"), ("1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1000", "0011", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0010", "0011", "0100", "0100", "0100", "0001", "0000", "0000", "0010", "0100", "1000", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "0111", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0010", "0010", "0011", "0011", "0001", "0001", "0000", "0000", "0010", "0111", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "0100", "0001", "0000", "0000", "0010", "0001", "0001", "0001", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "0101", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "0011", "0001", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0011", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0000", "0000", "0001", "0001", "0010", "0001", "0000", "0000", "0001", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0000", "0000", "0010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0000", "0000", "0001", "0001", "0010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0001", "0001", "0000", "0000", "0010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "1001"), ("1001", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0011", "0001", "0000", "0001", "0001", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0001", "0001", "0000", "0000", "0011", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "1000"), ("1001", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "0100", "0001", "0000", "0001", "0001", "0010", "0011", "0001", "0000", "0000", "0000", "0000", "0001", "0011", "0001", "0001", "0000", "0000", "0000", "0101", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1001", "0111", "0001", "0000", "0000", "0001", "0001", "0010", "0011", "0010", "0001", "0001", "0010", "0011", "0010", "0001", "0001", "0000", "0000", "0000", "1000", "1001", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1010", "0011", "0000", "0000", "0001", "0001", "0001", "0010", "0010", "0011", "0011", "0010", "0010", "0001", "0001", "0000", "0000", "0000", "0011", "1010", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1001", "1000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "1000", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000"), ("1000", "0111", "0111", "1001", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1010", "0101", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0001", "0110", "1010", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "1000", "1001", "0111", "0111", "1000"), ("1000", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1010", "0101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0101", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0110", "0111", "1000"), ("1000", "1000", "0111", "0110", "0110", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1010", "0111", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0111", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "1000", "1000"), ("1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1010", "1010", "0111", "0100", "0010", "0001", "0001", "0010", "0100", "0111", "1010", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001"), ("1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001"), ("0011", "0011", "0011", "0011", "0010", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0110", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0110", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0010", "0010", "0011", "0011", "0011"), ("0011", "0011", "0011", "0000", "0001", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0101", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0001", "0000", "0011", "0011", "0011"), ("0011", "0011", "0010", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0000", "0000", "0010", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "0000", "0000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0010", "0011", "0011"), ("0011", "0011", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0011", "0011"), ("0011", "0011", "0011", "0010", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0000", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0010", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"), ("0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011"));	 
begin


	--CIRCUIT 1: CONTROL GENERATOR
	--Static signals for DAC:
	 BLANKn <= '1'; --no blanking
	 SYNCn <= '0'; --no sync on green
	 --Create VGA clock (50MHz -> 25MHz):
	 process (clk)
	 begin
		 if rising_edge(clk) then
			clk_vga <= not clk_vga;
		 end if;
	 end process;
	 
	 --Create horizontal signals:
	 process (clk_vga)
		variable Hcount: natural range 0 to H_LOW + HBP + H_HIGH + HFP;
	begin
	 if rising_edge(clk_vga) then
		 Hcount := Hcount + 1;
		 if Hcount = H_LOW then
			Hsyn <= '1';
		 elsif Hcount = H_LOW + HBP then
			Hactive <= '1';
		 elsif Hcount = H_LOW + HBP + H_HIGH then
			Hactive <= '0';
		 elsif Hcount = H_LOW + HBP + H_HIGH + HFP then
			Hsyn <= '0';
			Hcount := 0;
		end if;
	end if;
end process;
 Hsync <= Hsyn; --internal signal converted to output

 
 --Create vertical signals:
 process (Hsyn)
	 variable Vcount: natural range 0 to V_LOW + VBP + V_HIGH + VFP;
 begin
	 if rising_edge(Hsyn) then
		Vcount := Vcount + 1;
		if Vcount = V_LOW then
			Vsyn <= '1';
		elsif Vcount = V_LOW + VBP then
			Vactive <= '1';
		elsif Vcount = V_LOW + VBP + V_HIGH then
			Vactive <= '0';
		elsif Vcount = V_LOW + VBP + V_HIGH + VFP then
			 Vsyn <= '0';
			 Vcount := 0;
		end if;
	 end if;
 end process;
 Vsync <= Vsyn; --not needed for Vsync; done just to match what was done to Hsync
 
 
 --Enable display:
 dena <= Hactive and Vactive;
 
 --CIRCUIT 2: IMAGE GENERATOR
 process (all)
	variable line_count: natural range 0 to V_HIGH;
	variable x: natural range 0 to H_HIGH;
	variable y: natural range 0 to V_HIGH;
	variable count: natural := 0;
 begin 
	 if rising_edge(Hsyn) then
		if Vactive then
			y := y + 1;
		 else
			y := 0;
		 end if;
	 end if;
	 if rising_edge(clk_vga) then
		if Hactive then
			x := x + 1;
		else
			x := 0;
		end if;
	 end if;
	 
	 if dena then
			if (y < 48 and x < 48) then
         R <= r_image_data(y)(x)(3 downto 0);
			G <= g_image_data(y)(x)(3 downto 0);
			B <= b_image_data(y)(x)(3 downto 0);
			else
			R <= (others => '0');
			 G <= (others => '0');
			 B <= (others => '0');
			end if;
			
		 else
			 R <= (others => '0');
			 G <= (others => '0');
			 B <= (others => '0');
		 end if;
	 end process;
end architecture;
---------------------

 

