//////////////////////////////////////////////////////////////////////
// Created by Actel SmartDesign Mon Jul 31 12:33:32 2023
// Testbench Template
// This is a basic testbench that instantiates your design with basic 
// clock and reset pins connected.  If your design has special
// clock/reset or testbench driver requirements then you should 
// copy this file and modify it. 
//////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps

module usr_testbench;

parameter SYSCLK_PERIOD = 22; // ~45MHz

reg SYSCLK;
reg NSYSRESET;
integer i;
reg [15:0] input_data;
wire [15:0] output_data;
initial
begin
    SYSCLK = 1'b0;
    NSYSRESET = 1'b1;
    input_data = 16'b0;
end

//////////////////////////////////////////////////////////////////////
// Reset Pulse
//////////////////////////////////////////////////////////////////////
initial
begin
    #(SYSCLK_PERIOD * 10 )
        NSYSRESET = 1'b0;
end


//////////////////////////////////////////////////////////////////////
// 10MHz Clock Driver
//////////////////////////////////////////////////////////////////////
always @(SYSCLK)
    #(SYSCLK_PERIOD / 2.0) SYSCLK <= !SYSCLK;


//////////////////////////////////////////////////////////////////////
// Instantiate Unit Under Test:  top
//////////////////////////////////////////////////////////////////////
peak_detection top_0 (
    // Inputs
    .input_data(input_data),
    .clk(SYSCLK),
    .reset(NSYSRESET),

    // Outputs
    .output_data(output_data)

    // Inouts

);
initial 
begin
    for (i=1; i < 20; i = i + 1)
    begin
        #(SYSCLK_PERIOD * 20)
            input_data = input_data + 1;
    end
    for (i=1; i < 20; i = i + 1)
    begin
        #(SYSCLK_PERIOD * 20)
            input_data = input_data - 1;
    end
	 for (i=1; i < 20; i = i + 1)
    begin
        #(SYSCLK_PERIOD * 20)
            input_data = input_data + 1;
	 end
	 for (i=1; i < 20; i = i + 1)
    begin
        #(SYSCLK_PERIOD * 20)
            input_data = input_data - 1;
	 end

end



endmodule

