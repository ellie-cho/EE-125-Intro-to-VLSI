module optiver (input [31:0] X, Y, output [31:0] Z);
assign Z = X ** 32;

endmodule